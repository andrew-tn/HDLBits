//https://hdlbits.01xz.net/wiki/Module_name

module top_module ( 
    input a, 
    input b, 
    input c,
    input d,
    output out1,
    output out2
);

endmodule
